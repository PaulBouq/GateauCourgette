//---------------------------------------------
// BE de l'UV 5.5 / 5.6 : Sécurisation d'un système SCADA
// Paul BOUQUET - Cédric DELAUNAY - Mathieu LOGARIO
//---------------------------------------------

//--------------------------------------------------
//                 Events
//--------------------------------------------------
event evt_send_ADMIN_WRITE_GC is        { send ADMIN_WRITE_GC from {env}1 to {GC}1 }
event evt_send_ADMIN_WRITE_LC1 is       { send ADMIN_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_ADMIN_WRITE_LC2 is       { send ADMIN_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_ADMIN_READ_GC is         { send ADMIN_READ_GC from {env}1 to {GC}1 }
event evt_send_ADMIN_READ_LC1 is        { send ADMIN_READ_LC1 from {env}1 to {GC}1 }
event evt_send_ADMIN_READ_LC2 is        { send ADMIN_READ_LC2 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_WRITE_GC is     { send GC_OWNER_WRITE_GC from {env}1 to {GC}1 }
event evt_send_GC_OWNER_WRITE_LC1 is    { send GC_OWNER_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_WRITE_LC2 is    { send GC_OWNER_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_READ_GC is      { send GC_OWNER_READ_GC from {env}1 to {GC}1 }
event evt_send_GC_OWNER_READ_LC1 is     { send GC_OWNER_READ_LC1 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_READ_LC2 is     { send GC_OWNER_READ_LC2 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_WRITE_GC is    { send LC1_OWNER_WRITE_GC from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_WRITE_LC1 is   { send LC1_OWNER_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_WRITE_LC2 is   { send LC1_OWNER_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_READ_GC is     { send LC1_OWNER_READ_GC from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_READ_LC1 is    { send LC1_OWNER_READ_LC1 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_READ_LC2 is    { send LC1_OWNER_READ_LC2 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_WRITE_GC is    { send LC2_OWNER_WRITE_GC from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_WRITE_LC1 is   { send LC2_OWNER_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_WRITE_LC2 is   { send LC2_OWNER_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_READ_GC is     { send LC2_OWNER_READ_GC from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_READ_LC1 is    { send LC2_OWNER_READ_LC1 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_READ_LC2 is    { send LC2_OWNER_READ_LC2 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_WRITE_GC is      { send UNKNOWN_WRITE_GC from {env}1 to {GC}1 }
event evt_send_UNKNOWN_WRITE_LC1 is     { send UNKNOWN_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_WRITE_LC2 is     { send UNKNOWN_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_READ_GC is       { send UNKNOWN_READ_GC from {env}1 to {GC}1 }
event evt_send_UNKNOWN_READ_LC1 is      { send UNKNOWN_READ_LC1 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_READ_LC2 is      { send UNKNOWN_READ_LC2 from {env}1 to {GC}1 }

event evt_recv_ADMIN_ACK_GC_WRITE is    { receive ACK_WRITE_GC_FOR_ADMIN from {GC}1 to {env}1 }
event evt_recv_ADMIN_ACK_GC_READ  is    { receive ACK_READ_GC_FOR_ADMIN from {GC}1 to {env}1 }

event evt_recv_ADMIN_NACK_GC_WRITE is   { receive NACK_WRITE_GC_FOR_ADMIN from {GC}1 to {env}1 }
event evt_recv_ADMIN_NACK_GC_READ  is   { receive NACK_READ_GC_FOR_ADMIN from {GC}1 to {env}1 }

event evt_recv_GC_OWNER_ACK_GC_READ is  { receive ACK_READ_GC_FOR_GC_OWNER from {GC}1 to {env}1 }

event evt_recv_LC1_OWNER_ACK_LC1_WRITE is {receive ACK_WRITE_LC1_FOR_LC1_OWNER from {GC}1 to {env}1 }
event evt_recv_LC1_OWNER_NACK_LC1_WRITE is {receive NACK_WRITE_LC1_FOR_LC1_OWNER from {GC}1 to {env}1 }
event evt_recv_LC2_OWNER_NACK_LC1_WRITE is {receive NACK_WRITE_LC1_FOR_LC2_OWNER from {GC}1 to {env}1 }

event evt_send_ADMIN_WRITE_NETWORK is {send ADMIN_WRITE_NETWORK from {env}1 to {GC}1 }
event evt_recv_ACK_WRITE_NETWORK_FROM_ADMIN is{receive ACK_WRITE_NETWORK_FROM_ADMIN from {GC}1 to {env}1 }


event evt_recv_LC1_OWNER_NACK_GC_READ is { receive NACK_READ_GC_FOR_LC1_OWNER from {GC}1 to {env}1 }
event evt_recv_LC2_OWNER_NACK_GC_READ is { receive NACK_READ_GC_FOR_LC2_OWNER from {GC}1 to {env}1 }
event evt_recv_UNKNOWN_NACK_GC_READ   is { receive NACK_READ_GC_FOR_UNKNOWN from {GC}1 to {env}1 }
event evt_recv_UNKNOWN_NACK_LC1_READ  is { receive NACK_READ_LC1_FOR_UNKNOWN from {GC}1 to {env}1 }
event evt_recv_UNKNOWN_NACK_LC2_READ  is { receive NACK_READ_LC2_FOR_UNKNOWN from {GC}1 to {env}1 }
event evt_recv_GC_OWNER_NACK_LC1_READ is { receive NACK_READ_LC1_FOR_GC_OWNER from {GC}1 to {env}1 }
event evt_recv_GC_OWNER_NACK_LC2_READ is { receive NACK_READ_LC1_FOR_GC_OWNER from {GC}1 to {env}1 }




event evt_recv_ANY is                   { receive ANY from {GC}1 to {env}1 }
event evt_send_END is                   { send REQ_END from {env}1 to {GC}1 }
event evt_recv_END is                   { receive REQ_END from {env}1 to {GC}1 }

//--------------------------------------------------
//           Activities Elementaires
//--------------------------------------------------

activity LC1_OWNER_READ_GC is
{
	event evt_send_LC1_OWNER_READ_GC; event evt_recv_LC1_OWNER_NACK_GC_READ
}

activity LC2_OWNER_READ_GC is
{
	event evt_send_LC2_OWNER_READ_GC; event evt_recv_LC2_OWNER_NACK_GC_READ
}

activity UNKNOWN_READ_GC is
{
	event evt_send_UNKNOWN_READ_GC; event evt_recv_UNKNOWN_NACK_GC_READ
}

activity UNKNOWN_READ_LC2 is
{
	event evt_send_UNKNOWN_READ_LC2; event evt_recv_UNKNOWN_NACK_LC2_READ
}

activity GC_OWNER_READ_LC1 is
{
	event evt_send_GC_OWNER_READ_LC1; event evt_recv_GC_OWNER_NACK_LC1_READ
}

activity GC_OWNER_READ_LC2 is
{
	event evt_send_GC_OWNER_READ_LC2; event evt_recv_GC_OWNER_NACK_LC2_READ
}


activity ADMIN_READ_GC is
{
    event evt_send_ADMIN_READ_GC; event evt_recv_ADMIN_ACK_GC_READ
}

activity GC_OWNER_READ_GC is
{
    event evt_send_GC_OWNER_READ_GC; event evt_recv_GC_OWNER_ACK_GC_READ
}

//--------------------------------------------------
//           Observateurs Elementaires
//--------------------------------------------------
property pty_actElem_ADMIN_WRITE_GC_allowed is 
{ 
  start   -- / / evt_send_ADMIN_WRITE_GC  /  -> waitRet;
  waitRet -- / / evt_recv_ADMIN_ACK_GC_WRITE  / -> start;
  waitRet -- / / evt_recv_ANY  /  -> reject
}

property pty_actElem_GC_OWNER_READ_GC_allowed is
{
    start -- / / evt_send_GC_OWNER_READ_GC / -> waitRet;
    waitRet -- / / evt_recv_GC_OWNER_ACK_GC_READ / -> start;
    waitRet -- / / evt_recv_ANY  /  -> reject
}

property pty_actElem_ADMIN_READ_GC_allowed is
{
    start -- / / evt_send_ADMIN_READ_GC / -> waitRet;
    waitRet -- / / evt_recv_ADMIN_ACK_GC_READ / -> start;
    waitRet -- / / evt_recv_ANY  /  -> reject
}

property pty_actElem_LC1OWNER_READ_GC_refused is
{
    start -- / / evt_send_LC1_OWNER_READ_GC / -> waitRet;
    waitRet -- / / evt_recv_LC1_OWNER_NACK_GC_READ / -> start;
    waitRet -- / / evt_recv_ANY / -> reject
}

property pty_actElem_LC2OWNER_READ_GC_refused is
{
    start -- / / evt_send_LC2_OWNER_READ_GC / -> waitRet;
    waitRet -- / / evt_recv_LC2_OWNER_NACK_GC_READ / -> start;
    waitRet -- / / evt_recv_ANY / -> reject
}

property pty_actElem_UNKNOWN_READ_GC_refused is
{
    start -- / / evt_send_UNKNOWN_READ_GC / -> waitRet;
    waitRet -- / / evt_recv_UNKNOWN_NACK_GC_READ / -> start;
    waitRet -- / / evt_recv_ANY / -> reject
}

//--------------------------------------------------
//              Contextes
//--------------------------------------------------

cdl confidentiality_Context_UNKNOWN_read_GC is
{
	properties
        pty_actElem_UNKNOWN_READ_GC_refused

	main is
	{
        UNKNOWN_READ_GC
    }
}

cdl confidentiality_Context_LC1OWNER_read_GC is
{
	properties
        pty_actElem_LC1OWNER_READ_GC_refused

	main is
	{
        LC1_OWNER_READ_GC
    }
}

cdl confidentiality_Context_LC2OWNER_read_GC is
{
	properties
        pty_actElem_LC2OWNER_READ_GC_refused

	main is
	{
        LC2_OWNER_READ_GC
    }
}


cdl availability_Context_ADMIN_read_GC is
{
    properties
        pty_actElem_ADMIN_READ_GC_allowed

    main is
    {
        ADMIN_READ_GC
    }
}

cdl availability_Context_GCOWNER_read_GC is
{
    properties
        pty_actElem_GC_OWNER_READ_GC_allowed        

    main is
    {
        GC_OWNER_READ_GC
    }
}