//---------------------------------------------
// BE de l'UV 5.5 / 5.6 : Sécurisation d'un système SCADA
// Paul BOUQUET - Cédric DELAUNAY - Mathieu LOGARIO
//---------------------------------------------

//--------------------------------------------------
//         Predicats 
//--------------------------------------------------

//--------------------------------------------------
//                 Events
//--------------------------------------------------
event evt_send_ADMIN_WRITE_GC is        { send ADMIN_WRITE_GC from {env}1 to {GC}1 }
event evt_send_ADMIN_WRITE_LC1 is       { send ADMIN_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_ADMIN_WRITE_LC2 is       { send ADMIN_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_ADMIN_READ_GC is         { send ADMIN_READ_GC from {env}1 to {GC}1 }
event evt_send_ADMIN_READ_LC1 is        { send ADMIN_READ_LC1 from {env}1 to {GC}1 }
event evt_send_ADMIN_READ_LC2 is        { send ADMIN_READ_LC2 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_WRITE_GC is     { send GC_OWNER_WRITE_GC from {env}1 to {GC}1 }
event evt_send_GC_OWNER_WRITE_LC1 is    { send GC_OWNER_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_WRITE_LC2 is    { send GC_OWNER_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_READ_GC is      { send GC_OWNER_READ_GC from {env}1 to {GC}1 }
event evt_send_GC_OWNER_READ_LC1 is     { send GC_OWNER_READ_LC1 from {env}1 to {GC}1 }
event evt_send_GC_OWNER_READ_LC2 is     { send GC_OWNER_READ_LC2 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_WRITE_GC is    { send LC1_OWNER_WRITE_GC from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_WRITE_LC1 is   { send LC1_OWNER_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_WRITE_LC2 is   { send LC1_OWNER_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_READ_GC is     { send LC1_OWNER_READ_GC from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_READ_LC1 is    { send LC1_OWNER_READ_LC1 from {env}1 to {GC}1 }
event evt_send_LC1_OWNER_READ_LC2 is    { send LC1_OWNER_READ_LC2 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_WRITE_GC is    { send LC2_OWNER_WRITE_GC from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_WRITE_LC1 is   { send LC2_OWNER_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_WRITE_LC2 is   { send LC2_OWNER_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_READ_GC is     { send LC2_OWNER_READ_GC from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_READ_LC1 is    { send LC2_OWNER_READ_LC1 from {env}1 to {GC}1 }
event evt_send_LC2_OWNER_READ_LC2 is    { send LC2_OWNER_READ_LC2 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_WRITE_GC is      { send UNKNOWN_WRITE_GC from {env}1 to {GC}1 }
event evt_send_UNKNOWN_WRITE_LC1 is     { send UNKNOWN_WRITE_LC1 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_WRITE_LC2 is     { send UNKNOWN_WRITE_LC2 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_READ_GC is       { send UNKNOWN_READ_GC from {env}1 to {GC}1 }
event evt_send_UNKNOWN_READ_LC1 is      { send UNKNOWN_READ_LC1 from {env}1 to {GC}1 }
event evt_send_UNKNOWN_READ_LC2 is      { send UNKNOWN_READ_LC2 from {env}1 to {GC}1 }

event evt_recv_ADMIN_ACK_GC_WRITE is    { receive ACK_WRITE_GC_FOR_ADMIN from {GC}1 to {env}1 }
event evt_recv_ADMIN_ACK_GC_READ  is    { receive ACK_READ_GC_FOR_ADMIN from {GC}1 to {env}1 }

event evt_recv_ADMIN_NACK_GC_WRITE is   { receive NACK_WRITE_GC_FOR_ADMIN from {GC}1 to {env}1 }
event evt_recv_ADMIN_NACK_GC_READ  is   { receive NACK_READ_GC_FOR_ADMIN from {GC}1 to {env}1 }


event evt_recv_ANY is                   { receive ANY from {GC}1 to {env}1 }
event evt_send_END is                   { send REQ_END from {env}1 to {GC}1 }
event evt_recv_END is                   { receive REQ_END from {env}1 to {GC}1 }

//--------------------------------------------------
//           Activities Elementaires
//--------------------------------------------------
activity actElem_ADMIN_WRITE_GC is 
{ event evt_send_ADMIN_WRITE_GC; { event evt_recv_ADMIN_ACK_GC_WRITE [] event evt_recv_ADMIN_NACK_GC_WRITE }
} 

//--------------------------------------------------
//           Observateurs Elementaires
//--------------------------------------------------
property pty_actElem_ADMIN_WRITE_GC_allowed is 
{ 
  start   -- / / evt_send_ADMIN_WRITE_GC  /  -> waitRet;
  waitRet -- / / evt_recv_ADMIN_ACK_GC_WRITE  / -> success;
  waitRet -- / / evt_recv_ANY  /  -> reject
}

//--------------------------------------------------
//              Contextes
//--------------------------------------------------
cdl cdl_my_Context is
{
    properties
        pty_actElem_ADMIN_WRITE_GC_allowed

    main is
    {
        actElem_ADMIN_WRITE_GC
    }
}